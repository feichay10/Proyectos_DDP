//Memoria de programa, se inicializa y no se modifica

module memprog(input  wire        clk,
               input  wire [9:0]  a,
               output wire [31:0] rd);

  reg [31:0] mem[0:1023]; //memoria de 1024 palabras de 32 bits de ancho

  initial
  begin
    $readmemb("//home//alumno//Escritorio//CPU_base//progfile.dat",mem); // inicializa la memoria del fichero en texto binario
  end
  
  assign rd = mem[a];

endmodule


